`include "packet.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "environment.sv"
