interface traffic_intf (input logic clock);
  
  
  logic reset;
  logic RED,GREEN,YELLOW;
endinterface

